`timescale 1ns / 1ps
//////////////////////////////////////////////////////////////////////////////////
// Company: 
// Engineer: Omar Ashraf Abd El Mongy
// 
// Create Date: 12/09/2024 08:56:08 PM
// Design Name: 
// Module Name: aes_ahb_interface
// Project Name: 
// Target Devices: 
// Tool Versions: 
// Description: 
// 
// Dependencies: 
// 
// Revision:
// Revision 0.01 - File Created
// Additional Comments:
// 
//////////////////////////////////////////////////////////////////////////////////
module aes_ahb_interface (
    input wire        HCLK,           // AHB Clock
    input wire        HRESETn,        // AHB Reset (active low)
    input wire        HSEL,           // AHB Select
    input wire [31:0] HADDR,          // AHB Address
    input wire        HWRITE,         // AHB Write Enable
    input wire        HREADY,         // AHB Ready
    input wire [31:0] HWDATA,         // AHB Write Data
    output reg [31:0] HRDATA,         // AHB Read Data
    output reg        HRESP,          // AHB Response
    input             DONE,           // AES Operation Done

    // Signals to AES Core
    output reg [127:0] aes_key,       // 128-bit Key
    output reg [127:0] aes_plaintext, // 128-bit Plaintext
    input  wire [127:0] aes_ciphertext,// 128-bit Ciphertext
    output reg         start          // Start Signal to AES Core
);
    // Address decoding for AES registers
    localparam KEY0_ADDR   = 32'h0000;
    localparam KEY1_ADDR   = 32'h0004;
    localparam KEY2_ADDR   = 32'h0008;
    localparam KEY3_ADDR   = 32'h000C;
    localparam TEXT0_ADDR  = 32'h0010;
    localparam TEXT1_ADDR  = 32'h0014;
    localparam TEXT2_ADDR  = 32'h0018;
    localparam TEXT3_ADDR  = 32'h001C;
    localparam CTRL_ADDR   = 32'h0020;
    localparam CIPHER0_ADDR = 32'h0024;
    localparam CIPHER1_ADDR = 32'h0028;
    localparam CIPHER2_ADDR = 32'h002C;
    localparam CIPHER3_ADDR = 32'h0030;

    reg [31:0] key_regs[3:0];        // 32-bit key registers
    reg [31:0] plaintext_regs[3:0]; // 32-bit plaintext registers

    // Register read/write logic
    always @(posedge HCLK or negedge HRESETn) begin
        HRESP <= DONE;
        if (!HRESETn) begin
            key_regs[0] <= 32'd0;
            key_regs[1] <= 32'd0;
            key_regs[2] <= 32'd0;
            key_regs[3] <= 32'd0;
            plaintext_regs[0] <= 32'd0;
            plaintext_regs[1] <= 32'd0;
            plaintext_regs[2] <= 32'd0;
            plaintext_regs[3] <= 32'd0;
            aes_key <= 128'd0;
            aes_plaintext <= 128'd0;
            HRDATA <= 32'd0;
            HRESP <= 1'b0;
            start <= 1'b0;
            //DONE <= 1'b0;
        end else if (HSEL && HREADY) begin
            if (HWRITE) begin
                // Write to registers
                case (HADDR)
                    KEY0_ADDR:  key_regs[0] <= HWDATA;
                    KEY1_ADDR:  key_regs[1] <= HWDATA;
                    KEY2_ADDR:  key_regs[2] <= HWDATA;
                    KEY3_ADDR:  key_regs[3] <= HWDATA;
                    TEXT0_ADDR: plaintext_regs[0] <= HWDATA;
                    TEXT1_ADDR: plaintext_regs[1] <= HWDATA;
                    TEXT2_ADDR: plaintext_regs[2] <= HWDATA;
                    TEXT3_ADDR: plaintext_regs[3] <= HWDATA;
                    CTRL_ADDR:  start <= HWDATA[0]; // Start encryption
                    default: ;
                endcase
            end else begin
                // Read from registers
                case (HADDR)
                    KEY0_ADDR:     HRDATA <= key_regs[0];
                    KEY1_ADDR:     HRDATA <= key_regs[1];
                    KEY2_ADDR:     HRDATA <= key_regs[2];
                    KEY3_ADDR:     HRDATA <= key_regs[3];
                    TEXT0_ADDR:    HRDATA <= plaintext_regs[0];
                    TEXT1_ADDR:    HRDATA <= plaintext_regs[1];
                    TEXT2_ADDR:    HRDATA <= plaintext_regs[2];
                    TEXT3_ADDR:    HRDATA <= plaintext_regs[3];
                    CIPHER0_ADDR:  HRDATA <= aes_ciphertext[31:0];
                    CIPHER1_ADDR:  HRDATA <= aes_ciphertext[63:32];
                    CIPHER2_ADDR:  HRDATA <= aes_ciphertext[95:64];
                    CIPHER3_ADDR:  HRDATA <= aes_ciphertext[127:96];
                    default:       HRDATA <= 32'd0;
                endcase
            end
        end
    end

    // Concatenate key and plaintext when all words are written
    always @(posedge HCLK or negedge HRESETn) begin
        if (!HRESETn) begin
            aes_key <= 128'd0;
            aes_plaintext <= 128'd0;
        end else begin
            aes_key <= {key_regs[3], key_regs[2], key_regs[1], key_regs[0]};
            aes_plaintext <= {plaintext_regs[3], plaintext_regs[2], plaintext_regs[1], plaintext_regs[0]};
        end
    end
endmodule

